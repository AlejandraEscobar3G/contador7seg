library verilog;
use verilog.vl_types.all;
entity contador7seg_vlg_vec_tst is
end contador7seg_vlg_vec_tst;
